--- !ruby/object:Hangman::Game
word: TERRAZZO
display_word: TERRA___
guessed_wrong:
- F
- H
- N
- Q
- S
num_wrong: 5
