--- !ruby/object:Hangman::Game
word: PARVE
display_word: ____E
guessed_wrong:
- S
num_wrong: 1
